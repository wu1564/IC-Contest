module geofence_v3 (  //with a modified booth multiplier
	clk,
	reset,
	X,
	Y,
	valid,
	is_inside
);

input clk;
input reset;
input [9:0] X;
input [9:0] Y;
output reg valid;
output reg is_inside;

////////////////////Parameters//////////////////////
localparam IDLE = 4'd0;
localparam RECEIVE = 4'd1;
localparam CREATE_VECTOR = 4'd2;
localparam CROSS_PRODUCT_STAGE_1 = 4'd3;
localparam CROSS_PRODUCT_STAGE_2 = 4'd4;
localparam JUDGE = 4'd5;
localparam TWO_VECTOR = 4'd6;
localparam CROSS_PRODUCT2_STAGE_1 = 4'd7;
localparam CROSS_PRODUCT2_STAGE_2 = 4'd8;
localparam JUDGE2 = 4'd9;
localparam FINAL = 4'd10;
////////////////////////////////////////////////////

//////////////Private Declaration///////////////////
// necessary
reg [9:0] target_x;
reg [9:0] target_y;
reg [9:0] point_x[0:5];
reg [9:0] point_y[0:5];
// my algorithm used 
wire start_flag_wire;
wire strobe;
wire signed [11:0] multiplicand_wire;
wire signed [11:0] multiplier_wire;
wire signed [23:0] result;
reg start_flag;
reg [3:0] state, next_state;
reg [2:0] receive_cnt, cycle_cnt;
reg [2:0] record;
reg signed [10:0] vector_x[0:1];
reg signed [10:0] vector_y[0:1];
reg signed [10:0] multiplicand;
reg signed [10:0] multiplier;
reg signed [21:0] calculate;
////////////////////////////////////////////////////

//*********************module***********************
modified_booth multiply(
	.clk(clk),
	.reset(reset),
	//.multiplicand({{1{multiplicand_wire[10]}},multiplicand_wire}),  // multiplicand * multiplier
	.multiplicand(multiplicand_wire),  // multiplicand * multiplier
	.multiplier(multiplier_wire),
	.result(result),
	.start_flag(start_flag_wire),
	.strobe(strobe)	
);
//**************************************************

///////////////////////wires////////////////////////
assign start_flag_wire = start_flag;
assign multiplicand_wire = {multiplicand[10],multiplicand};
assign multiplier_wire = {multiplier[10],multiplier};
////////////////////////////////////////////////////

////////////////////start_flag//////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		start_flag <= 1'b0;
	end else begin
		case (state) 
			CROSS_PRODUCT_STAGE_1, 
			CROSS_PRODUCT_STAGE_2, 
			CROSS_PRODUCT2_STAGE_1, 
			CROSS_PRODUCT2_STAGE_2: start_flag <= (receive_cnt == 3'd0) ? 1'b1 : 1'b0;
	    	default: 				start_flag <= 1'b0;
		endcase
	end
end
////////////////////////////////////////////////////

/////////////////multiplicand///////////////////////	
always @(posedge clk or posedge reset) begin
	if(reset) begin
		multiplicand <= 11'd0;
	end else begin
		case (state)             // vec_x[0] * vec_y[1] - vec_x[1] * vec_y[0]
			CROSS_PRODUCT_STAGE_1, CROSS_PRODUCT2_STAGE_1:  multiplicand <= vector_x[0];
			CROSS_PRODUCT_STAGE_2, CROSS_PRODUCT2_STAGE_2:  multiplicand <= vector_x[1];
	    	default: multiplicand <= multiplicand;
		endcase
	end
end
////////////////////////////////////////////////////

//////////////////////multiplier////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		multiplier <= 11'd0;
	end else begin
		case (state)             // vec_x[0] * vec_y[1] - vec_x[1] * vec_y[0]
			CROSS_PRODUCT_STAGE_1, CROSS_PRODUCT2_STAGE_1:  multiplier <= vector_y[1];
			CROSS_PRODUCT_STAGE_2, CROSS_PRODUCT2_STAGE_2:  multiplier <= vector_y[0];
	    	default: multiplier <= multiplier;
		endcase
	end
end
////////////////////////////////////////////////////

//////////////////////next_state////////////////////
always @(*) begin
	case (state) 
	    IDLE: 					next_state = RECEIVE;
	    RECEIVE:				next_state = (receive_cnt == 3'd5) ? CREATE_VECTOR : RECEIVE;
	    CREATE_VECTOR: 			next_state = (record != 3'd4) ? CROSS_PRODUCT_STAGE_1 : TWO_VECTOR;
	    CROSS_PRODUCT_STAGE_1:	next_state = (strobe) ? CROSS_PRODUCT_STAGE_2 : CROSS_PRODUCT_STAGE_1;
	    CROSS_PRODUCT_STAGE_2: 	next_state = (strobe) ? JUDGE : CROSS_PRODUCT_STAGE_2;
	    JUDGE:					next_state = CREATE_VECTOR;
	    TWO_VECTOR:				next_state = (cycle_cnt == 3'd6) ? FINAL : CROSS_PRODUCT2_STAGE_1;
	    CROSS_PRODUCT2_STAGE_1: next_state = (strobe) ? CROSS_PRODUCT2_STAGE_2 : CROSS_PRODUCT2_STAGE_1;
	    CROSS_PRODUCT2_STAGE_2: next_state = (strobe) ? JUDGE2 : CROSS_PRODUCT2_STAGE_2;
	    JUDGE2:					next_state = TWO_VECTOR;
	    FINAL:					next_state = (cycle_cnt == 3'd1) ? IDLE : FINAL;
	    default:				next_state = IDLE;
	endcase
end
////////////////////////////////////////////////////

//////////////////////state/////////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		state <= IDLE;
	end else begin
		state <= next_state;
	end
end
////////////////////////////////////////////////////

//////////////////////receive_cnt///////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		receive_cnt <= 3'd0;
	end else begin
		case (state)
			RECEIVE: 				receive_cnt <= receive_cnt + 3'd1;
			CROSS_PRODUCT_STAGE_1,
			CROSS_PRODUCT_STAGE_2,
			CROSS_PRODUCT2_STAGE_1,
			CROSS_PRODUCT2_STAGE_2: receive_cnt <= (strobe) ? 3'd0 : 3'd1;
			default: 				receive_cnt <= 3'd0;
		endcase
	end
end
////////////////////////////////////////////////////

///////////////////////target_x/////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		target_x <= 10'd0;
	end else begin
		case (state)
			IDLE: 	 target_x <= X;
			default: target_x <= target_x; 
		endcase
	end
end
////////////////////////////////////////////////////

///////////////////////target_y/////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		target_y <= 10'd0;
	end else begin
		case (state)
			IDLE:	 target_y <= Y;
			default: target_y <= target_y;
		endcase
	end
end
////////////////////////////////////////////////////

//////////////////////point_x///////////////////////
integer i;
always @(posedge clk or posedge reset) begin
	if(reset) begin
		for(i = 0; i < 6; i = i + 1) begin
			point_x[i] <= 10'd0;
		end
	end else begin
		case (state)
			RECEIVE:	point_x[receive_cnt] <= X;
			JUDGE:		begin
							if(~calculate[21]) begin
								case (cycle_cnt) 
									3'd0:		begin
													point_x[1] <= point_x[2];
													point_x[2] <= point_x[1];
												end
									3'd1:		begin
													point_x[2] <= point_x[3];
													point_x[3] <= point_x[2];
												end
									3'd2:		begin
													point_x[3] <= point_x[4];
													point_x[4] <= point_x[3];
												end			
									3'd3:		begin
													point_x[4] <= point_x[5];
													point_x[5] <= point_x[4];
												end
								    default:	begin
													for(i = 0; i < 6; i = i + 1) begin
														point_x[i] <= point_x[i];
													end
								    			end
								endcase
							end
						end
			default:	begin
							for(i = 0; i < 6; i = i + 1) begin
								point_x[i] <= point_x[i];
							end
						end
		endcase
	end
end
////////////////////////////////////////////////////

//////////////////////point_y///////////////////////
integer j;
always @(posedge clk or posedge reset) begin
	if(reset) begin
		for(j = 0; j < 6; j = j + 1) begin
			point_y[j] <= 10'd0;
		end
	end else begin
		case (state)
			RECEIVE:	point_y[receive_cnt] <= Y;
			JUDGE:		begin
							if(~calculate[21]) begin
								case (cycle_cnt) 
									3'd0:		begin
													point_y[1] <= point_y[2];
													point_y[2] <= point_y[1];
												end
									3'd1:		begin
													point_y[2] <= point_y[3];
													point_y[3] <= point_y[2];
												end
									3'd2:		begin
													point_y[3] <= point_y[4];
													point_y[4] <= point_y[3];
												end			
									3'd3:		begin
													point_y[4] <= point_y[5];
													point_y[5] <= point_y[4];
												end
								    default:	begin
								    				for(j = 0; j < 6; j = j + 1) begin
								    					point_y[j] <= point_y[j];
								    				end
								    			end
								endcase
							end
						end
			default:	begin
							for(j = 0; j < 6; j = j + 1) begin
								point_y[j] <= point_y[j];
							end
						end
		endcase
	end
end
////////////////////////////////////////////////////

///////////////////record/////////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		record <= 3'd0;
	end else begin
		case (state)
			IDLE:	 		record <= 3'd0;
			CREATE_VECTOR:	record <= (record == 3'd4) ? 3'd0 : record;
			JUDGE:	 		record <= (calculate[21]) ? record + 3'd1 : 3'd0;
			JUDGE2:			record <= (~calculate[21]) ? record + 3'd1 : record;
			default: 		record <= record;
		endcase
	end
end
////////////////////////////////////////////////////

/////////////////////cycle_cnt//////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		cycle_cnt <= 3'd0;
	end else begin
		case (state)
			IDLE:	 		cycle_cnt <= 3'd0;
			CREATE_VECTOR:	cycle_cnt <= (record == 3'd4) ? 3'd0 : cycle_cnt;
			JUDGE:	 		cycle_cnt <= (cycle_cnt != 3'd3) ? cycle_cnt + 3'd1 : 3'd0;
			JUDGE2:			cycle_cnt <= (cycle_cnt != 3'd6) ? cycle_cnt + 3'd1 : 3'd0;
			FINAL:			cycle_cnt <= 3'd1;
			default: 		cycle_cnt <= cycle_cnt;
		endcase
	end
end
////////////////////////////////////////////////////

////////////////////////vector_x////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		vector_x[0] <= 11'd0;
		vector_x[1] <= 11'd0;
	end else begin
		case (state) 
			CREATE_VECTOR: 	begin
								case (cycle_cnt) 
									3'd0:		begin
													vector_x[0] <= {1'b0,point_x[1]} - {1'b0,point_x[0]};
													vector_x[1] <= {1'b0,point_x[2]} - {1'b0,point_x[0]};			
												end
									3'd1:		begin
													vector_x[0] <= {1'b0,point_x[2]} - {1'b0,point_x[0]};
													vector_x[1] <= {1'b0,point_x[3]} - {1'b0,point_x[0]};			
												end
									3'd2:		begin
													vector_x[0] <= {1'b0,point_x[3]} - {1'b0,point_x[0]};
													vector_x[1] <= {1'b0,point_x[4]} - {1'b0,point_x[0]};			
												end
									3'd3:		begin
													vector_x[0] <= {1'b0,point_x[4]} - {1'b0,point_x[0]};
													vector_x[1] <= {1'b0,point_x[5]} - {1'b0,point_x[0]};			
												end
								    default:	begin
								    				vector_x[0] <= vector_x[0];
								    				vector_x[1] <= vector_x[1];
								    			end
								endcase
							end
			TWO_VECTOR:		begin
								case (cycle_cnt)
									3'd0:		begin
													vector_x[0] <= {1'b0,target_x} - {1'b0,point_x[0]};
													vector_x[1] <= {1'b0,point_x[1]} - {1'b0,point_x[0]};			
												end
									3'd1:		begin
													vector_x[0] <= {1'b0,target_x} - {1'b0,point_x[1]};
													vector_x[1] <= {1'b0,point_x[2]} - {1'b0,point_x[1]};			
												end
									3'd2:		begin
													vector_x[0] <= {1'b0,target_x} - {1'b0,point_x[2]};
													vector_x[1] <= {1'b0,point_x[3]} - {1'b0,point_x[2]};			
												end
									3'd3:		begin
													vector_x[0] <= {1'b0,target_x} - {1'b0,point_x[3]};
													vector_x[1] <= {1'b0,point_x[4]} - {1'b0,point_x[3]};			
												end
									3'd4:		begin
													vector_x[0] <= {1'b0,target_x} - {1'b0,point_x[4]};
													vector_x[1] <= {1'b0,point_x[5]} - {1'b0,point_x[4]};			
												end
									3'd5:		begin
													vector_x[0] <= {1'b0,target_x} - {1'b0,point_x[5]};
													vector_x[1] <= {1'b0,point_x[0]} - {1'b0,point_x[5]};
												end
									default:	begin
													vector_x[0] <= vector_x[0];
													vector_x[1] <= vector_x[1];
												end
								endcase
							end
		    default: 		begin
		    					vector_x[0] <= vector_x[0];
		    					vector_x[1] <= vector_x[1];	
		    				end
		endcase
	end
end
////////////////////////////////////////////////////

////////////////////////vector_y////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		vector_y[0] <= 11'd0;
		vector_y[1] <= 11'd0;
	end else begin
		case (state) 
			CREATE_VECTOR: 	begin
								vector_y[0] <= {1'b0,point_y[cycle_cnt + 3'd1]} - {1'b0,point_y[0]};
								vector_y[1] <= {1'b0,point_y[cycle_cnt + 3'd2]} - {1'b0,point_y[0]};		
							end
			TWO_VECTOR:		begin
								case (cycle_cnt)
									3'd5:		begin
													vector_y[0] <= {1'b0,target_y} - {1'b0,point_y[5]};
													vector_y[1] <= {1'b0,point_y[0]} - {1'b0,point_y[5]};
												end
									3'd6:		begin
													vector_y[0] <= vector_y[0];
													vector_y[1] <= vector_y[1];
												end
									default:	begin
													vector_y[0] <= {1'b0,target_y} - {1'b0,point_y[cycle_cnt]};
													vector_y[1] <= {1'b0,point_y[cycle_cnt + 3'd1]} - {1'b0,point_y[cycle_cnt]};			
												end
								endcase
							end
		    default: 		begin
		    					vector_y[0] <= vector_y[0];
		    					vector_y[1] <= vector_y[1];	
		    				end
		endcase
	end
end
////////////////////////////////////////////////////

///////////////////////calculate////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		calculate <= 22'd0;
	end else begin
		case (state)       //vec_x[0] * vec_y[1] - vec_x[1] * vec_y[0]
			CROSS_PRODUCT_STAGE_1, CROSS_PRODUCT2_STAGE_1:	calculate <= result[21:0];
			CROSS_PRODUCT_STAGE_2, CROSS_PRODUCT2_STAGE_2:	calculate <= (strobe) ? calculate - result[21:0] : calculate;
		    default: calculate <= calculate;
		endcase
	end
end
////////////////////////////////////////////////////

///////////////////////valid////////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		valid <= 1'b0;
	end else begin
		case (state)
			FINAL: 	 valid <= (cycle_cnt == 3'd1) ? 1'b0 : 1'b1;
			default: valid <= 1'b0;
		endcase
	end
end
///////////////////////////////////////////////////////

/////////////////////is_inside/////////////////////////
always @(posedge clk or posedge reset) begin
	if(reset) begin
		is_inside <= 1'b0;
	end else begin
		case (state) 
			FINAL:	 is_inside <= (cycle_cnt != 3'd1) ? (record == 3'd6) ? 1'b1 : 1'b0 : 1'd0;
		    default: is_inside <= 1'b0;
		endcase
	end
end
////////////////////////////////////////////////////

endmodule
